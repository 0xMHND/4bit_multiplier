*** SPICE deck for cell 4bit_multiplier{sch} from library Multiplier
*** Created on Mon Mar 13, 2017 23:39:41
*** Last revised on Fri Mar 17, 2017 19:05:13
*** Written on Fri Mar 17, 2017 19:05:40 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS



*** SUBCIRCUIT Gates_v2__nand2-bb_2-sz_10 FROM CELL Gates_v2:nand2{sch}
.SUBCKT Gates_v2__nand2-bb_2-sz_10 A A_NAND_B B
** GLOBAL gnd
** GLOBAL vdd
XNMOS@0 A_NAND_B B net@64 NMOS W='WW*4*(1+ABN/sqrt(WW*4*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*4*(Lwid))'
XNMOS@1 net@64 A gnd NMOS W='WW*4*(1+ABN/sqrt(WW*4*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*4*(Lwid))'
XPMOS@0 A_NAND_B B vdd  PMOS W='WW*5*(1+ABN/sqrt(WW*5*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*5*(Lwid))'
XPMOS@1 A_NAND_B A vdd  PMOS W='WW*5*(1+ABN/sqrt(WW*5*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*5*(Lwid))'
.ENDS Gates_v2__nand2-bb_2-sz_10

*** SUBCIRCUIT Gates_v2__xor2 FROM CELL Gates_v2:xor2{sch}
.SUBCKT Gates_v2__xor2 A A_NAND_B A_XOR_B B
** GLOBAL gnd
** GLOBAL vdd
Xnand2@9 A net@12 A_NAND_B Gates_v2__nand2-bb_2-sz_10
Xnand2@10 net@75 A_XOR_B net@12 Gates_v2__nand2-bb_2-sz_10
Xnand2@11 A_NAND_B net@75 B Gates_v2__nand2-bb_2-sz_10
Xnand2@12 A A_NAND_B B Gates_v2__nand2-bb_2-sz_10
.ENDS Gates_v2__xor2

*** SUBCIRCUIT Adder__1bit_adder_v2 FROM CELL Adder:1bit_adder_v2{sch}
.SUBCKT Adder__1bit_adder_v2 A B Cin Cout sum
** GLOBAL gnd
** GLOBAL vdd
Xnand2@0 net@13 Cout net@15 Gates_v2__nand2-bb_2-sz_10
Xxor2@0 A net@15 net@4 B Gates_v2__xor2
Xxor2@1 net@4 net@13 sum Cin Gates_v2__xor2
.ENDS Adder__1bit_adder_v2

*** SUBCIRCUIT Adder__4bit_adder FROM CELL Adder:4bit_adder{sch}
.SUBCKT Adder__4bit_adder A0 A1 A2 A3 B0 B1 B2 B3 Cin Cout sum0 sum1 sum2 sum3
** GLOBAL gnd
** GLOBAL vdd
X_1bit_add@0 A0 B0 Cin net@7 sum0 Adder__1bit_adder_v2
X_1bit_add@5 A1 B1 net@7 net@41 sum1 Adder__1bit_adder_v2
X_1bit_add@8 A2 B2 net@41 net@46 sum2 Adder__1bit_adder_v2
X_1bit_add@9 A3 B3 net@46 Cout sum3 Adder__1bit_adder_v2
.ENDS Adder__4bit_adder

*** SUBCIRCUIT Gates_v2__nand3-bb_2-sz_10 FROM CELL Gates_v2:nand3{sch}
.SUBCKT Gates_v2__nand3-bb_2-sz_10 A A_AND_B_AND_C B C gnd vdd
** GLOBAL gnd
** GLOBAL vdd
XNMOS@0 A_AND_B_AND_C A net@2 NMOS W='WW*4*(1+ABN/sqrt(WW*4*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*4*(Lwid))'
XNMOS@1 net@2 B net@22 NMOS W='WW*4*(1+ABN/sqrt(WW*4*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*4*(Lwid))'
XNMOS@2 net@22 C gnd NMOS W='WW*4*(1+ABN/sqrt(WW*4*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*4*(Lwid))'
XPMOS@0 A_AND_B_AND_C A vdd  PMOS W='WW*4*(1+ABN/sqrt(WW*4*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*4*(Lwid))'
XPMOS@1 A_AND_B_AND_C B vdd  PMOS W='WW*4*(1+ABN/sqrt(WW*4*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*4*(Lwid))'
XPMOS@2 A_AND_B_AND_C C vdd  PMOS W='WW*4*(1+ABN/sqrt(WW*4*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*4*(Lwid))'
.ENDS Gates_v2__nand3-bb_2-sz_10

*** SUBCIRCUIT Multiplier__D_flipflop FROM CELL Multiplier:D_flipflop{sch}
.SUBCKT Multiplier__D_flipflop clk Data Q _Q
** GLOBAL gnd
** GLOBAL vdd
Xnand2@1 clk net@5 net@0 Gates_v2__nand2-bb_2-sz_10
Xnand2@2 net@5 net@0 net@12 Gates_v2__nand2-bb_2-sz_10
Xnand2@5 Data net@12 net@42 Gates_v2__nand2-bb_2-sz_10
Xnand2@6 net@42 _Q Q Gates_v2__nand2-bb_2-sz_10
Xnand2@7 _Q Q net@5 Gates_v2__nand2-bb_2-sz_10
Xnand3@0 net@5 net@42 clk net@12 gnd vdd Gates_v2__nand3-bb_2-sz_10
.ENDS Multiplier__D_flipflop

*** SUBCIRCUIT Multiplier__16bit-flipflop FROM CELL Multiplier:16bit-flipflop{sch}
.SUBCKT Multiplier__16bit-flipflop clk d0 d1 d10 d11 d12 d13 d14 d15 d2 d3 d4 d5 d6 d7 d8 d9 q0 q1 q10 q11 q12 q13 q14 q15 q2 q3 q4 q5 q6 q7 q8 q9
** GLOBAL gnd
** GLOBAL vdd
XD_flipfl@0 clk d2 q2 D_flipfl@0__Q Multiplier__D_flipflop
XD_flipfl@1 clk d1 q1 D_flipfl@1__Q Multiplier__D_flipflop
XD_flipfl@2 clk d0 q0 D_flipfl@2__Q Multiplier__D_flipflop
XD_flipfl@3 clk d3 q3 D_flipfl@3__Q Multiplier__D_flipflop
XD_flipfl@4 clk d6 q6 D_flipfl@4__Q Multiplier__D_flipflop
XD_flipfl@5 clk d5 q5 D_flipfl@5__Q Multiplier__D_flipflop
XD_flipfl@6 clk d4 q4 D_flipfl@6__Q Multiplier__D_flipflop
XD_flipfl@7 clk d7 q7 D_flipfl@7__Q Multiplier__D_flipflop
XD_flipfl@8 clk d10 q10 D_flipfl@8__Q Multiplier__D_flipflop
XD_flipfl@9 clk d9 q9 D_flipfl@9__Q Multiplier__D_flipflop
XD_flipfl@10 clk d8 q8 D_flipfl@10__Q Multiplier__D_flipflop
XD_flipfl@11 clk d11 q11 D_flipfl@11__Q Multiplier__D_flipflop
XD_flipfl@12 clk d14 q14 D_flipfl@12__Q Multiplier__D_flipflop
XD_flipfl@13 clk d13 q13 D_flipfl@13__Q Multiplier__D_flipflop
XD_flipfl@14 clk d12 q12 D_flipfl@14__Q Multiplier__D_flipflop
XD_flipfl@15 clk d15 q15 D_flipfl@15__Q Multiplier__D_flipflop
.ENDS Multiplier__16bit-flipflop

*** SUBCIRCUIT Gates_v2__inv-bb_2-sz_10 FROM CELL Gates_v2:inv{sch}
.SUBCKT Gates_v2__inv-bb_2-sz_10 gnd in out vdd
** GLOBAL gnd
** GLOBAL vdd
XNMOS@0 out in gnd NMOS W='WW*3*(1+ABN/sqrt(WW*3*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*3*(Lwid))'
XPMOS@0 out in vdd  PMOS W='WW*6.667*(1+ABN/sqrt(WW*6.667*(Lwid)))' L='(Lwid)' DELVTO='AVT0N/sqrt(WW*6.667*(Lwid))'
.ENDS Gates_v2__inv-bb_2-sz_10

*** SUBCIRCUIT Gates_v2__and2 FROM CELL Gates_v2:and2{sch}
.SUBCKT Gates_v2__and2 A A_AND_B B
** GLOBAL gnd
** GLOBAL vdd
Xinv@0 gnd net@0 A_AND_B vdd Gates_v2__inv-bb_2-sz_10
Xnand2@0 A net@0 B Gates_v2__nand2-bb_2-sz_10
.ENDS Gates_v2__and2

.global gnd vdd

*** SUBCIRCUIT _4bit_multiplier FROM CELL Multiplier:4bit_multiplier{sch}
.SUBCKT _4bit_multiplier A0 A1 A2 A3 B0 B1 B2 B3 Cin clk gnd sum0 sum1 sum2 sum3 sum4 sum5 sum6 sum7
** GLOBAL gnd
** GLOBAL vdd
X_4bit_add@0 net@558 net@559 net@560 net@561 net@73 net@144 net@75 net@139 Cin net@566 net@562 net@563 net@564 net@565 Adder__4bit_adder
X_4bit_add@2 net@555 net@556 net@557 gnd net@29 net@30 net@31 net@32 Cin net@534 net@587 net@530 net@531 net@588 Adder__4bit_adder
X_4bit_add@3 net@567 net@570 net@568 net@569 net@103 net@152 net@105 net@153 Cin sum7 sum3 sum4 sum5 sum6 Adder__4bit_adder
X_16bit-fl@0 clk A0 A1 gnd gnd B0 B1 B2 B3 A2 A3 gnd gnd gnd gnd gnd gnd net@336 net@340 _16bit-fl@0_q10 _16bit-fl@0_q11 net@298 net@299 net@471 net@466 net@344 net@348 _16bit-fl@0_q4 _16bit-fl@0_q5 _16bit-fl@0_q6 _16bit-fl@0_q7 _16bit-fl@0_q8 _16bit-fl@0_q9 Multiplier__16bit-flipflop
X_16bit-fl@1 clk net@336 net@340 gnd gnd gnd gnd net@471 net@466 net@344 net@348 net@467 net@587 net@530 net@531 net@588 net@534 net@408 net@412 _16bit-fl@1_q10 _16bit-fl@1_q11 _16bit-fl@1_q12 _16bit-fl@1_q13 net@399 net@465 net@416 net@420 net@485 net@490 net@558 net@559 net@560 net@561 Multiplier__16bit-flipflop
X_16bit-fl@2 clk net@408 net@412 net@566 gnd gnd gnd gnd net@465 net@416 net@420 net@485 net@490 net@562 net@563 net@564 net@565 A0 A1 net@569 _16bit-fl@2_q11 _16bit-fl@2_q12 _16bit-fl@2_q13 _16bit-fl@2_q14 net@116 A2 A3 sum0 sum1 sum2 net@567 net@570 net@568 Multiplier__16bit-flipflop
Xand2@0 net@336 net@467 net@298 Gates_v2__and2
Xand2@1 net@340 net@555 net@298 Gates_v2__and2
Xand2@2 net@344 net@556 net@298 Gates_v2__and2
Xand2@3 net@348 net@557 net@298 Gates_v2__and2
Xand2@4 net@336 net@29 net@299 Gates_v2__and2
Xand2@5 net@340 net@30 net@299 Gates_v2__and2
Xand2@6 net@344 net@31 net@299 Gates_v2__and2
Xand2@7 net@348 net@32 net@299 Gates_v2__and2
Xand2@8 net@408 net@73 net@399 Gates_v2__and2
Xand2@9 net@412 net@144 net@399 Gates_v2__and2
Xand2@10 net@416 net@75 net@399 Gates_v2__and2
Xand2@11 net@420 net@139 net@399 Gates_v2__and2
Xand2@16 A0 net@103 net@116 Gates_v2__and2
Xand2@17 A1 net@152 net@116 Gates_v2__and2
Xand2@18 A2 net@105 net@116 Gates_v2__and2
Xand2@19 A3 net@153 net@116 Gates_v2__and2
.ENDS _4bit_multiplier


X_4bit_multiplier A0 A1 A2 A3 B0 B1 B2 B3 Cin clk gnd sum0 sum1 sum2 sum3 sum4 sum5 sum6 sum7 _4bit_multiplier

.END
