*** SPICE deck for cell 4bit_adder{sch} from library Adder
*** Created on Tue Feb 28, 2017 18:27:12
*** Last revised on Thu Mar 02, 2017 18:48:45
*** Written on Thu Mar 02, 2017 18:54:44 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS

*** SUBCIRCUIT Gates_v2__nand2 FROM CELL Gates_v2:nand2{sch}
.SUBCKT Gates_v2__nand2 A A_NAND_B B
** GLOBAL gnd
** GLOBAL vdd
XNMOS@0 A_NAND_B B net@64 NMOS
XNMOS@1 net@64 A gnd NMOS
XPMOS@0 A_NAND_B B vdd PMOS
XPMOS@1 A_NAND_B A vdd PMOS
.ENDS Gates_v2__nand2

*** SUBCIRCUIT Gates_v2__xor2 FROM CELL Gates_v2:xor2{sch}
.SUBCKT Gates_v2__xor2 A A_NAND_B A_XOR_B B
** GLOBAL gnd
** GLOBAL vdd
Xnand2@9 A net@12 A_NAND_B Gates_v2__nand2
Xnand2@10 net@75 A_XOR_B net@12 Gates_v2__nand2
Xnand2@11 A_NAND_B net@75 B Gates_v2__nand2
Xnand2@12 A A_NAND_B B Gates_v2__nand2
.ENDS Gates_v2__xor2

*** SUBCIRCUIT Adder__1bit_adder_v2 FROM CELL 1bit_adder_v2{sch}
.SUBCKT Adder__1bit_adder_v2 A B Cin Cout sum
** GLOBAL gnd
** GLOBAL vdd
Xnand2@0 net@13 Cout net@15 Gates_v2__nand2
Xxor2@0 A net@15 net@4 B Gates_v2__xor2
Xxor2@1 net@4 net@13 sum Cin Gates_v2__xor2
.ENDS Adder__1bit_adder_v2

.global gnd vdd

*** TOP LEVEL CELL: 4bit_adder{sch}
X_1bit_add@0 A0 B0 Cin net@7 sum0 Adder__1bit_adder_v2
X_1bit_add@5 A1 B1 net@7 net@41 sum1 Adder__1bit_adder_v2
X_1bit_add@8 A2 B2 net@41 net@46 sum2 Adder__1bit_adder_v2
X_1bit_add@9 A3 B3 net@46 Cout sum3 Adder__1bit_adder_v2
.END
